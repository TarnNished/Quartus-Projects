module xor_gate(z,x,y);
input x,y;
output z;
xor (z,x,y);
endmodule